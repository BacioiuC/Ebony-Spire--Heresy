return {
-- Table: {1}
{
   ["soundVolume"]=-0.11,
   ["fullScreen"]=false,
   ["uiZoomToggle"]=false,
},
}